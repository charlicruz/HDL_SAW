--------------------------------------------------------------------------------
-- Company: 
-- Engineer:
--
-- Create Date:   12:43:04 07/15/2020
-- Design Name:   
-- Module Name:   Y:/carlos ITEFI/ITEFI-PROYECTOS/HDL_SAW/MOJO/genera_clock/test.vhd
-- Project Name:  genera
-- Target Device:  
-- Tool versions:  
-- Description:   
-- 
-- VHDL Test Bench Created by ISE for module: PWM_COUNTER
-- 
-- Dependencies:
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
--
-- Notes: 
-- This testbench has been automatically generated using types std_logic and
-- std_logic_vector for the ports of the unit under test.  Xilinx recommends
-- that these types always be used for the top-level I/O of a design in order
-- to guarantee that the testbench will bind correctly to the post-implementation 
-- simulation model.
--------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
 
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--USE ieee.numeric_std.ALL;
 
ENTITY test IS
END test;
 
ARCHITECTURE behavior OF test IS 
 
    -- Component Declaration for the Unit Under Test (UUT)
 
    COMPONENT PWM_COUNTER
    PORT(
         CLK : IN  std_logic;
         RST : IN  std_logic;
         PWM_IN : IN  std_logic;
         PWM_COUNT : OUT  std_logic_vector(15 downto 0)
        );
    END COMPONENT;
    

   --Inputs
   signal CLK : std_logic := '0';
   signal RST : std_logic := '0';
   signal PWM_IN : std_logic := '0';

 	--Outputs
   signal PWM_COUNT : std_logic_vector(15 downto 0);

   -- Clock period definitions
   constant CLK_period : time := 10 ns;
 
BEGIN
 
	-- Instantiate the Unit Under Test (UUT)
   uut: PWM_COUNTER PORT MAP (
          CLK => CLK,
          RST => RST,
          PWM_IN => PWM_IN,
          PWM_COUNT => PWM_COUNT
        );

   -- Clock process definitions
   CLK_process :process
   begin
		CLK <= '0';
		wait for CLK_period/2;
		CLK <= '1';
		wait for CLK_period/2;
   end process;
 

   -- Stimulus process
   stim_proc: process
   begin		
      -- hold reset state for 100 ns.
      wait for 100 ns;	

      wait for CLK_period*10;
     
      -- insert stimulus here 
      PWM_IN <= '0';
		wait for CLK_period*10;
		PWM_IN <= '1';
		wait for CLK_period*10;
		PWM_IN <= '0';
--		wait for CLK_period*4;
--		PWM_IN <= '1';
--		wait for CLK_period*4;
--		PWM_IN <= '0';
--		wait for CLK_period*4;
--		PWM_IN <= '1';
--		wait for CLK_period*4;
--      wait;
   end process;

END;
