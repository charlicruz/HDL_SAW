--library ieee;
--use ieee.std_logic_1164.all;
--use ieee.std_logic_arith.all;
--use ieee.std_logic_unsigned.all;
--use ieee.numeric_std.all;
--use work.myPaquete.all;
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.std_logic_unsigned.all;
use ieee.std_logic_arith.all;

entity ssgdemo is
	Port (	entrada : in std_logic;
	         mclk	:	in		std_logic;
			--	led0	:	out	std_logic;
				pwm0		:	out	std_logic;
				pwm1		:	out	std_logic;
				pwm2		:	out	std_logic;
				pwm3		:	out	std_logic;
				pwm4		:	out	std_logic;
				pwm5		:	out	std_logic;                                                                                                                                                                                              
			--	seleccion_mux : in std_logic_vector(7 down to 0);
				reset : in std_logic;
				aux_coun : out STD_LOGIC_VECTOR (3 downto 0);--std_logic;
				data_difference : out STD_LOGIC_VECTOR (3 downto 0);--std_logic;
--				cntr2	:	out		std_logic_vector (1 downto 0);
				aux_coun2 : out STD_LOGIC_VECTOR (3 downto 0);--std_logic;
				data_difference2 : out STD_LOGIC_VECTOR (3 downto 0);--std_logic;
			--	mclkout :	out	std_logic;
			--	cclkout:	out	std_logic;
				clk,rst : in  STD_LOGIC;
			   led : out  STD_LOGIC_VECTOR (7 downto 0);
				dec : out  STD_LOGIC_VECTOR (4 downto 0);
	--		   spi_ss,spi_mosi,spi_sck,avr_tx,avr_rx_busy : in STD_LOGIC;
				rx    : in std_logic;
				tx : out std_logic;
				--sigdel: out std_logic;
--				sigdel:IN std_logic;
--			   entrada_xor:IN std_logic;
		--		seleccion_mux: in std_logic_vector (1 downto 0);
				signal2: out std_logic;
			   salida: out  STD_LOGIC_VECTOR (7 downto 0)

				);
end ssgdemo;

architecture Behaivioral of ssgdemo is
signal clkdiv	:		std_logic_vector(28 downto 0);
signal cntr0	:		std_logic_vector(6 downto 0);
signal cntr1	:		std_logic_vector(6 downto 0);
signal cntr2	:		std_logic_vector(6 downto 0);
signal cntr3	:		std_logic_vector(6 downto 0);--nuevo
signal cntrv	:		std_logic_vector(6 downto 0);
signal pwmclk	:		std_logic;
signal cclk		:		std_logic;
signal cntclk	:		std_logic;
--signal cclkout	:		std_logic;
--signal mclkout	:		std_logic;
signal seleccion_mux : std_logic_vector (2 downto 0):=(others=>'0');
signal cnt 		: 		UNSIGNED(6 downto 0);
signal pwmv		:		std_logic;
signal contador : STD_LOGIC_VECTOR (26 downto 0) :=B"000000000000000000000000000";  --Hex 50M=2FAF080
--signal leds     : STD_LOGIC_VECTOR (7 downto  0) :=B"00000000";

signal aux_count : STD_LOGIC_VECTOR (3 downto  0) :=B"0000";--std_logic;-- := '0';
signal entrada_xor : std_logic := '0';	
signal sigDel : std_logic:= '0';
signal count_xor : STD_LOGIC_VECTOR (3 downto  0):=B"0000";--std_logic;
signal aux_count2 : STD_LOGIC_VECTOR (3 downto  0) :=B"0000";--std_logic;-- := '0';
signal entrada_xor2 : std_logic := '0';	
signal sigDel2 : std_logic:= '0';
signal count_xor2 : STD_LOGIC_VECTOR (3 downto  0);--:=B"0000";--std_logic;

signal digit    : std_logic;
signal segments : STD_LOGIC_VECTOR (7 downto  0);--:=B"0000";--std_logic;


signal auxiliar1    : std_logic;
signal predeterminado1    : std_logic;


signal clk_18432_s : std_logic                    := '0';
signal data_s      : std_logic_vector(7 downto 0) := x"00";
signal in_valid_s  : std_logic                    := '0';
signal out_valid_s : std_logic                    := '0';
signal accept_s    : std_logic                    := '0';
signal tx_s : std_logic                    := '0';
signal rx_s    : std_logic                    := '0';	
signal temporal: STD_LOGIC;
signal temporal2: STD_LOGIC;
signal temporal3: STD_LOGIC;

signal conta: integer range 0 to 124999 := 0;
signal mux_out: STD_LOGIC;
signal salidaff1: STD_LOGIC;--_vector (3 downto 0);
signal salidaff2: STD_LOGIC;
signal salidaff3: STD_LOGIC;
signal salidaff4: STD_LOGIC;
signal salidaff5: STD_LOGIC;
signal salidaff6: STD_LOGIC;
signal salidaff7: STD_LOGIC;

signal b:std_logic_vector(3 downto 0);
signal p:std_logic_vector(4 downto 0); 
component CLKMIX is
port
 (-- Clock in ports
  CLK_IN1           : in     std_logic;
  -- Clock out ports
  CLK_OUT1          : out    std_logic
 );
end component;  

component clk_18432 is
port 
 (clk   : in std_logic;
  reset : in std_logic;
  clk_18432 : out std_logic);
end component clk_18432;

    component uart_tx is
        port (clk      : in std_logic;
              reset    : in std_logic;
              data_in  : in std_logic_vector(7 downto 0);
              in_valid : in std_logic;

              tx        : out std_logic;
              accept_in : out std_logic);
    end component uart_tx;

    component uart_rx is
        port (clk   : in std_logic;
              reset : in std_logic;
              rx    : in std_logic;

              data_out  : out std_logic_vector(7 downto 0);
              out_valid : out std_logic);
    end component uart_rx;


begin
  u1: CLKMIX port map
   (-- Clock in ports
    CLK_IN1 => mclk,
    -- Clock out ports
    CLK_OUT1 => cclk);
	 
	process (cclk)
			begin
				if cclk='1' and cclk'event then
					clkdiv <= clkdiv + 1;
				end if;
	end process;
	
	
--	cclkout <= cclk;
--	mclkout <= mclk;

	pwmclk <= clkdiv(4);
	cntclk <= clkdiv (24);
--	led0   <= clkdiv(10);
	

--	se�al1: process(clk,rst)
--	begin
--		if rising_edge(clk) then
--			if (rst='1') then
--				auxiliar1 <= '0';
--				aux_count <= (others=>'0');
--			elsif rising_edge(entrada) then
--				if (contador=124999) then
--				auxiliar1 <= not(temporal1);
--				aux_count <= 0);
--			else
--				aux_count <= aux_count+'1';
--			end if;
--		end if;
--	end process;
--		
--	se�al1: process(clk,rst,aux_count)
--	begin
--		if rising_edge(clk) then
--			if (rst='1') then
--				auxiliar1 <= '0';
--				aux_count <= (others=>'0');
--			elsif (aux_count=predeterminado1) then
--				auxiliar1 <= not auxiliar1;
--				aux_count <= (others=>'0');
--			else
--				aux_count <= aux_count+'1';
--			end if;
--		end if;
--	end process;
	
	process (cntclk)
			begin
			if cntclk = '1' and cntclk'event then -- duty
						cntr0 <= cntr0 + 1;
						cntrv <= cntrv + 1;
						cntr1 <= "0000001";
						cntr2 <= "0000001";
						cntr3 <= "0000010";
				end if;
		end process;
	
	 process (rst, entrada) begin
        if (rst = '1') then
            temporal <= '0';
				 temporal2 <= '0';
            conta <= 0;
        elsif rising_edge(entrada) then
            if (conta = 124) then--124999
                temporal <= NOT(temporal);
					 temporal2 <= temporal after 1200ns;
					 temporal3 <= temporal after 1800ns;
                conta <= 0;
            else
                conta <= conta+1;
            end if;
        end if;
    end process;
  
--    process (rst, entrada) begin
--        if (rst = '1') then
--            temporal2 <= '0';
--            conta <= 0;
--        elsif rising_edge(entrada) then
--            if (conta = 120) then--124999
--                temporal2 <= NOT(temporal2);
--                conta <= 0;
--            else
--                conta <= conta+1;
--            end if;
--        end if;
--    end process;    
	 pwm5<=temporal;
    pwm4 <= temporal2;
	 pwm3<=temporal3;
	 process(seleccion_mux,temporal,salidaff1,salidaff2,salidaff3,salidaff4,salidaff5,salidaff6,salidaff7)
	 begin
		case seleccion_mux is
			when "000" => mux_out<=temporal;
			when "001" => mux_out<=salidaff1;
			when "010" => mux_out<=salidaff2;
			when "011" => mux_out<=salidaff3;
			when "100" => mux_out<=salidaff4;
			when "101" => mux_out<='0';--salidaff5;
			when "110" => mux_out<=salidaff6; 
			when "111" => mux_out<=salidaff7;
			when others=> mux_out<='0';
		end case;
	 end process;
	 --pwm3<=mux_out;
	 
	process(pwmclk, reset) begin
        if reset = '0' then
            cnt <= (others => '0');
        elsif rising_edge(pwmclk) then
            if cnt = 99 then --99 then -- 320MHz /2 = 160MHz / 99 = 1.62MHz
               -- temporal <= NOT(temporal);
					 cnt <= (others => '0');				 
            else
                cnt <= cnt + 1;
            end if;
        end if;
    end process;
		
	 pwmv <= '1' when (cnt < UNSIGNED(cntrv)) else '0';
	 pwm0 <= '1' when (cnt < UNSIGNED(cntr0)) else '0';
	 pwm1 <= '1' when (cnt < UNSIGNED(cntr1)) else '0';
	-- pwm3 <= '1' when (cnt < UNSIGNED(cntr3)) else '0';
		
	process(pwmv) begin
		if pwmv = '0' and cnt < UNSIGNED(cntr2) then
			pwm2 <= '1';			
		else
			pwm2 <= '0';
		
		end if;
	end process;
	
	data_difference <= count_xor;
   data_difference2 <= count_xor2;
	entrada_xor2<=temporal3 xor temporal;
	entrada_xor<=temporal2 xor temporal;--temporal2;
	sigDel<=temporal;
	contador_xor:process(clk,entrada_xor,sigDel)
		begin
			if falling_edge(clk) then
				if entrada_xor='1' then
					aux_count<= aux_count+1;
				elsif ( entrada_xor='0' and sigDel='1') then
					count_xor<=aux_count;
					aux_count<=(others=>'0');
				end if;
				if entrada_xor2='1' then
					aux_count2<= aux_count2+1;
				elsif ( entrada_xor2='0' and sigDel2='1') then
					count_xor2<=aux_count2;
					aux_count2<=(others=>'0');
				end if;
			sigDel<=entrada_xor;
			sigDel2<=entrada_xor2;

			end if;
	end process;
   aux_coun<= aux_count;
	aux_coun2<= aux_count2;

b<=aux_count;

binbcd4:process(b,p)
begin
p(4)<= (b(3) and b(2)) or (b(3) and b(1));
p(3)<= (b(3) and not b(2) and not b(1)); 
p(2)<= (not b(3) and b(2)) or (b(2) and b(1)); 
p(1)<= (b(3) and b(2) and not b(1)) or (not b(3) and b(1));-- and b(1));
p(0)<= b(0);
end process;
dec<=p;

 process(p)
	 begin
		case p is
			when "00000" => segments<="11000000";
			when "00001" => segments<="11111001";
			when "00010" => segments<="10100100";
			when "00011" => segments<="10110000";
			when "00100" => segments<="11000000";
			when "00101" => segments<="10011001";
			when "00110" => segments<="10010010"; 
			when "00111" => segments<="10000011";
			when "01000" => segments<="11111000";
			when "01001" => segments<="10011000";
			when others  => segments<="11111111";
		end case;
	 end process;
--tx<=segments;
in_valid_s <= accept_s and out_valid_s;
    
    clk_gen : clk_18432 port map (clk   => clk,
                                  reset => reset,

                                  clk_18432 => clk_18432_s);

    tx_0 : uart_tx port map (clk      => clk_18432_s,
                             reset    => reset,
                             data_in  => data_s,
                             in_valid => in_valid_s,

                             tx        => tx,
                             accept_in => accept_s);

    rx_0 : uart_rx port map (clk   => clk_18432_s,
                             reset => reset,
                             rx    => rx,

                             data_out  => data_s,
                             out_valid => out_valid_s); 
end Behaivioral;
		